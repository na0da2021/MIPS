module adder( input  [31:0] data_in1, data_in2,
              output [31:0] result);

assign result = data_in1 + data_in2;
				  
endmodule